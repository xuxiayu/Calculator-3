package top_pkg;
   import uvm_pkg::*;
   
`include "env.sv"
`include "tests.sv"
endpackage // top_pkg
   