package top_pkg;

   import uvm_pkg::*;

   // include the env
   `include "env.sv"   
   
   // Define the sequences and tests 
   `include "tests.sv" 
   
endpackage // top_pkg
